    ����          Assembly-CSharp   Saves+Position   xyz      ףп{�>����